`timescale  1ns / 1ps

module InstructionMem (
         Address,
         dout
       );
input [8: 0] Address;
output [31: 0] dout;

	parameter MEM_SIZE = 512;
	reg [31:0]RAM[0:MEM_SIZE-1];
	
	assign dout = RAM[Address];

initial	begin
RAM[9'd0] <=  32'h 3c011001;
RAM[9'd1] <=  32'h 343a0000;
RAM[9'd2] <=  32'h 8f510000;
RAM[9'd3] <=  32'h 8f520004;
RAM[9'd4] <=  32'h 8f530008;
RAM[9'd5] <=  32'h 8f54000c;
RAM[9'd6] <=  32'h 001af025;
RAM[9'd7] <=  32'h 00006025;
RAM[9'd8] <=  32'h 0c100072;
RAM[9'd9] <=  32'h 218c0004;
RAM[9'd10] <=  32'h 200d0028;
RAM[9'd11] <=  32'h 0c10007c;
RAM[9'd12] <=  32'h 0c1000b6;
RAM[9'd13] <=  32'h 0c100099;
RAM[9'd14] <=  32'h 0c100072;
RAM[9'd15] <=  32'h 218c0004;
RAM[9'd16] <=  32'h 15acfffa;
RAM[9'd17] <=  32'h 0c10007c;
RAM[9'd18] <=  32'h 0c1000b6;
RAM[9'd19] <=  32'h 0c100072;
RAM[9'd20] <=  32'h 1000ffff;
RAM[9'd21] <=  32'h 01404825;
RAM[9'd22] <=  32'h 00002825;
RAM[9'd23] <=  32'h 20060004;
RAM[9'd24] <=  32'h 340400ff;
RAM[9'd25] <=  32'h 31210003;
RAM[9'd26] <=  32'h 312200fc;
RAM[9'd27] <=  32'h 005a1020;
RAM[9'd28] <=  32'h 8c420020;
RAM[9'd29] <=  32'h 00001825;
RAM[9'd30] <=  32'h 10610006;
RAM[9'd31] <=  32'h 20630001;
RAM[9'd32] <=  32'h 10610008;
RAM[9'd33] <=  32'h 20630001;
RAM[9'd34] <=  32'h 1061000a;
RAM[9'd35] <=  32'h 00441024;
RAM[9'd36] <=  32'h 08100030;
RAM[9'd37] <=  32'h 00042600;
RAM[9'd38] <=  32'h 00441024;
RAM[9'd39] <=  32'h 00021602;
RAM[9'd40] <=  32'h 08100030;
RAM[9'd41] <=  32'h 00042400;
RAM[9'd42] <=  32'h 00441024;
RAM[9'd43] <=  32'h 00021402;
RAM[9'd44] <=  32'h 08100030;
RAM[9'd45] <=  32'h 00042200;
RAM[9'd46] <=  32'h 00441024;
RAM[9'd47] <=  32'h 00021202;
RAM[9'd48] <=  32'h 2004ff00;
RAM[9'd49] <=  32'h 01645824;
RAM[9'd50] <=  32'h 01625825;
RAM[9'd51] <=  32'h 20a50001;
RAM[9'd52] <=  32'h 000b3a02;
RAM[9'd53] <=  32'h 000b4600;
RAM[9'd54] <=  32'h 00e85825;
RAM[9'd55] <=  32'h 00094a02;
RAM[9'd56] <=  32'h 14c5ffde;
RAM[9'd57] <=  32'h 03e00008;
RAM[9'd58] <=  32'h 100c0010;
RAM[9'd59] <=  32'h 00180a00;
RAM[9'd60] <=  32'h 00181602;
RAM[9'd61] <=  32'h 00225025;
RAM[9'd62] <=  32'h afdf02d8;
RAM[9'd63] <=  32'h 23de0004;
RAM[9'd64] <=  32'h 0c100015;
RAM[9'd65] <=  32'h 23defffc;
RAM[9'd66] <=  32'h 8fdf02d8;
RAM[9'd67] <=  32'h 019a7020;
RAM[9'd68] <=  32'h 8dc1011c;
RAM[9'd69] <=  32'h 01610826;
RAM[9'd70] <=  32'h 02a1a826;
RAM[9'd71] <=  32'h 02d5b026;
RAM[9'd72] <=  32'h 02f6b826;
RAM[9'd73] <=  32'h 0317c026;
RAM[9'd74] <=  32'h 03e00008;
RAM[9'd75] <=  32'h 8f550010;
RAM[9'd76] <=  32'h 8f560014;
RAM[9'd77] <=  32'h 8f570018;
RAM[9'd78] <=  32'h 8f58001c;
RAM[9'd79] <=  32'h 03e00008;
RAM[9'd80] <=  32'h 00c00825;
RAM[9'd81] <=  32'h 00003824;
RAM[9'd82] <=  32'h 00005024;
RAM[9'd83] <=  32'h 340b0004;
RAM[9'd84] <=  32'h 302200ff;
RAM[9'd85] <=  32'h 3023ff00;
RAM[9'd86] <=  32'h 00031a02;
RAM[9'd87] <=  32'h 00431026;
RAM[9'd88] <=  32'h 3c0300ff;
RAM[9'd89] <=  32'h 00231824;
RAM[9'd90] <=  32'h 00032c02;
RAM[9'd91] <=  32'h 00031bc2;
RAM[9'd92] <=  32'h 306400ff;
RAM[9'd93] <=  32'h 14640008;
RAM[9'd94] <=  32'h 00651826;
RAM[9'd95] <=  32'h 00431026;
RAM[9'd96] <=  32'h 3c03ff00;
RAM[9'd97] <=  32'h 00231824;
RAM[9'd98] <=  32'h 00031dc2;
RAM[9'd99] <=  32'h 306400ff;
RAM[9'd100] <=  32'h 14640003;
RAM[9'd101] <=  32'h 08100069;
RAM[9'd102] <=  32'h 3883001b;
RAM[9'd103] <=  32'h 0810005e;
RAM[9'd104] <=  32'h 3883001b;
RAM[9'd105] <=  32'h 00431026;
RAM[9'd106] <=  32'h 214a0001;
RAM[9'd107] <=  32'h 00073a00;
RAM[9'd108] <=  32'h 00e23825;
RAM[9'd109] <=  32'h 00014200;
RAM[9'd110] <=  32'h 00014e02;
RAM[9'd111] <=  32'h 01090825;
RAM[9'd112] <=  32'h 156affe3;
RAM[9'd113] <=  32'h 03e00008;
RAM[9'd114] <=  32'h afdf02d8;
RAM[9'd115] <=  32'h 23de0004;
RAM[9'd116] <=  32'h 0c10003a;
RAM[9'd117] <=  32'h 23defffc;
RAM[9'd118] <=  32'h 8fdf02d8;
RAM[9'd119] <=  32'h 02358826;
RAM[9'd120] <=  32'h 02569026;
RAM[9'd121] <=  32'h 02779826;
RAM[9'd122] <=  32'h 0298a026;
RAM[9'd123] <=  32'h 03e00008;
RAM[9'd124] <=  32'h 00115025;
RAM[9'd125] <=  32'h afdf02d8;
RAM[9'd126] <=  32'h 23de0004;
RAM[9'd127] <=  32'h 0c100015;
RAM[9'd128] <=  32'h 23defffc;
RAM[9'd129] <=  32'h 8fdf02d8;
RAM[9'd130] <=  32'h 000b8825;
RAM[9'd131] <=  32'h 00125025;
RAM[9'd132] <=  32'h afdf02d8;
RAM[9'd133] <=  32'h 23de0004;
RAM[9'd134] <=  32'h 0c100015;
RAM[9'd135] <=  32'h 23defffc;
RAM[9'd136] <=  32'h 8fdf02d8;
RAM[9'd137] <=  32'h 000b9025;
RAM[9'd138] <=  32'h 00135025;
RAM[9'd139] <=  32'h afdf02d8;
RAM[9'd140] <=  32'h 23de0004;
RAM[9'd141] <=  32'h 0c100015;
RAM[9'd142] <=  32'h 23defffc;
RAM[9'd143] <=  32'h 8fdf02d8;
RAM[9'd144] <=  32'h 000b9825;
RAM[9'd145] <=  32'h 00145025;
RAM[9'd146] <=  32'h afdf02d8;
RAM[9'd147] <=  32'h 23de0004;
RAM[9'd148] <=  32'h 0c100015;
RAM[9'd149] <=  32'h 23defffc;
RAM[9'd150] <=  32'h 8fdf02d8;
RAM[9'd151] <=  32'h 000ba025;
RAM[9'd152] <=  32'h 03e00008;
RAM[9'd153] <=  32'h 00113025;
RAM[9'd154] <=  32'h afdf02d8;
RAM[9'd155] <=  32'h 23de0004;
RAM[9'd156] <=  32'h 0c100050;
RAM[9'd157] <=  32'h 23defffc;
RAM[9'd158] <=  32'h 8fdf02d8;
RAM[9'd159] <=  32'h 00078825;
RAM[9'd160] <=  32'h 00123025;
RAM[9'd161] <=  32'h afdf02d8;
RAM[9'd162] <=  32'h 23de0004;
RAM[9'd163] <=  32'h 0c100050;
RAM[9'd164] <=  32'h 23defffc;
RAM[9'd165] <=  32'h 8fdf02d8;
RAM[9'd166] <=  32'h 00079025;
RAM[9'd167] <=  32'h 00133025;
RAM[9'd168] <=  32'h afdf02d8;
RAM[9'd169] <=  32'h 23de0004;
RAM[9'd170] <=  32'h 0c100050;
RAM[9'd171] <=  32'h 23defffc;
RAM[9'd172] <=  32'h 8fdf02d8;
RAM[9'd173] <=  32'h 00079825;
RAM[9'd174] <=  32'h 00143025;
RAM[9'd175] <=  32'h afdf02d8;
RAM[9'd176] <=  32'h 23de0004;
RAM[9'd177] <=  32'h 0c100050;
RAM[9'd178] <=  32'h 23defffc;
RAM[9'd179] <=  32'h 8fdf02d8;
RAM[9'd180] <=  32'h 0007a025;
RAM[9'd181] <=  32'h 03e00008;
RAM[9'd182] <=  32'h 3c0600ff;
RAM[9'd183] <=  32'h 3c07ff00;
RAM[9'd184] <=  32'h 34e7ffff;
RAM[9'd185] <=  32'h 3408ff00;
RAM[9'd186] <=  32'h 3c09ffff;
RAM[9'd187] <=  32'h 352900ff;
RAM[9'd188] <=  32'h 340a00ff;
RAM[9'd189] <=  32'h 3c0bffff;
RAM[9'd190] <=  32'h 356bff00;
RAM[9'd191] <=  32'h 02462824;
RAM[9'd192] <=  32'h 02270824;
RAM[9'd193] <=  32'h 00250825;
RAM[9'd194] <=  32'h 02682824;
RAM[9'd195] <=  32'h 00290824;
RAM[9'd196] <=  32'h 00250825;
RAM[9'd197] <=  32'h 028a2824;
RAM[9'd198] <=  32'h 002b0824;
RAM[9'd199] <=  32'h 00250825;
RAM[9'd200] <=  32'h 02662824;
RAM[9'd201] <=  32'h 02471024;
RAM[9'd202] <=  32'h 00451025;
RAM[9'd203] <=  32'h 02882824;
RAM[9'd204] <=  32'h 00491024;
RAM[9'd205] <=  32'h 00451025;
RAM[9'd206] <=  32'h 022a2824;
RAM[9'd207] <=  32'h 004b1024;
RAM[9'd208] <=  32'h 00451025;
RAM[9'd209] <=  32'h 02862824;
RAM[9'd210] <=  32'h 02671824;
RAM[9'd211] <=  32'h 00651825;
RAM[9'd212] <=  32'h 02282824;
RAM[9'd213] <=  32'h 00691824;
RAM[9'd214] <=  32'h 00651825;
RAM[9'd215] <=  32'h 024a2824;
RAM[9'd216] <=  32'h 006b1824;
RAM[9'd217] <=  32'h 00651825;
RAM[9'd218] <=  32'h 02262824;
RAM[9'd219] <=  32'h 02872024;
RAM[9'd220] <=  32'h 00852025;
RAM[9'd221] <=  32'h 02482824;
RAM[9'd222] <=  32'h 00892024;
RAM[9'd223] <=  32'h 00852025;
RAM[9'd224] <=  32'h 026a2824;
RAM[9'd225] <=  32'h 008b2024;
RAM[9'd226] <=  32'h 00852025;
RAM[9'd227] <=  32'h 00208825;
RAM[9'd228] <=  32'h 00409025;
RAM[9'd229] <=  32'h 00609825;
RAM[9'd230] <=  32'h 0080a025;
RAM[9'd231] <=  32'h 03e00008;


	end

endmodule
